module alu1(
    output result,
    output carryout,
    output zero,
    input A,
    input B,
    input carryin,
    input[7:0] command
)
