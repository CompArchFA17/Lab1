module mux2to1
(
  output      selected,
  input[1:0]  inputs,
  input       select
);

endmodule

module mux8to1
(
  output selected,
  input[7:0] inputs,
  input[2:0] select
);

endmodule