//Single bit slice module for ALU

module BitSlice(
    output cout, sum, res,
    input ADD, SUB, XOR, AND, NAND, NOR, OR, A, B, CIN
);
   

endmodule
