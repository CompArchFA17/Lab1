//Single bit slice module for ALU

module BitSlice
(
    output cout, sum, res,
    input ADD, SUB, XOR, AND, NAND, NOR, OR, A, B, CIN
);
    // TODO This is fake testing code
        assign cout = 0;
        assign res = 0;
        assign sum = 0;

endmodule
