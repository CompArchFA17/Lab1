// Implementation of an ALU that performs addition, subtraction, XOR, SLT, OR, NOR, NAND, and AND operations.

`include "operations.v"

// Definine command numbers
`define CADD  3'd0
`define CSUB  3'd1
`define CXOR  3'd2
`define CSLT  3'd3
`define CAND  3'd4
`define CNAND 3'd5
`define CNOR  3'd6
`define COR   3'd7

// Implementation of a control logic LUT to determine ALU operation.
module ALUcontrolLUT
(
output reg[2:0] 	muxindex,
output reg	invertB,
output reg	othercontrolsignal,
input[2:0]	ALUcommand
);

  always @(ALUcommand) begin
    case (ALUcommand)
      `CADD:  begin muxindex = 0; invertB=0; othercontrolsignal = 0; end
      `CSUB:  begin muxindex = 0; invertB=1; othercontrolsignal = 0; end
      `CXOR:  begin muxindex = 1; invertB=0; othercontrolsignal = 0; end
      `CSLT:  begin muxindex = 2; invertB=0; othercontrolsignal = 0; end
      `CAND:  begin muxindex = 3; invertB=0; othercontrolsignal = 0; end
      `CNAND: begin muxindex = 3; invertB=0; othercontrolsignal = 1; end
      `CNOR:  begin muxindex = 4; invertB=0; othercontrolsignal = 1; end
      `COR:   begin muxindex = 4; invertB=0; othercontrolsignal = 0; end
    endcase
  end
endmodule

// Define macros for second LUT.
`define MADDSUB 3'd0
`define MXOR 3'd1
`define MSLT 3'd2
`define MANDNAND 3'd3
`define MNOROR 3'd4

// Decide which operation results to output based on the results of the index 
// generated by the control LUT.
module ALUoutputLUT
(
input[31:0] operandA,
input[31:0] operandB,
input[2:0] muxindex,
input invertB,
input othercontrolsignal,
output reg[31:0] result,
output reg carryout,
output reg zero,
output reg overflow
);

// The results of each module.
wire[31:0] resAddsub;
wire[31:0] resXor;
wire[31:0] resSlt;
wire[31:0] resAndnand;
wire[31:0] resNoror;

// The carryout flags of each module.
wire carryoutAddSub;
wire carryoutXor;
wire carryoutSLT;
wire carryoutAND;
wire carryoutOR;

// The zero flags of each module.
wire zeroAddSub;
wire zeroXor;
wire zeroSLT;
wire zeroAND;
wire zeroOR;

// The overflow flags of each module.
wire overflowAddSub;
wire overflowXor;
wire overflowSLT;
wire overflowAND;
wire overflowOR;

AddSub #1000 dut0 (resAddsub, carryoutAddSub, zeroAddSub, overflowAddSub, operandA, operandB, invertB);
alu32bitxor dut1 (resXor, carryoutXor, zeroXor, overflowXor, operandA, operandB);
alu32bitslt dut2 (resSlt, carryoutSLT, zeroSLT, overflowSLT, operandA, operandB);
alu32bitandn dut3 (resAndnand, carryoutAND, zeroAND, overflowAND, operandA, operandB, othercontrolsignal);
NOROR dut4 (resNoror, carryoutOR, zeroOR, overflowOR, operandA, operandB, othercontrolsignal);

// The LUT behaves as a set of muxes that choose each bit of the result and each flag based on the muxindex 
// it is passed as an address.
always @(muxindex or resAddsub or resXor or resSlt or resAndnand or resNoror) begin
 case(muxindex)
    `MADDSUB: begin  result = resAddsub;   carryout = carryoutAddSub;  zero = zeroAddSub;  overflow = overflowAddSub; end
    `MXOR: begin     result = resXor;      carryout = carryoutXor;     zero = zeroXor;     overflow = overflowXor; end
    `MSLT: begin     result = resSlt;      carryout = carryoutSLT;     zero = zeroSLT;     overflow = overflowSLT; end
    `MANDNAND: begin result = resAndnand;  carryout = carryoutAND;     zero = zeroAND;     overflow = overflowAND; end
    `MNOROR: begin   result = resNoror;    carryout = carryoutOR;      zero = zeroOR;      overflow = overflowOR; end
  endcase
end

endmodule

// Implementation of the ALU in it's entirety.
module ALU
(
output[31:0]  result,
output        carryout,
output        zero,
output        overflow,
input[31:0]   operandA,
input[31:0]   operandB,
input[2:0]    command
);

wire[2:0]   muxindex;
wire  invertB;
wire othercontrolsignal;

ALUcontrolLUT controlLookup (muxindex, invertB, othercontrolsignal, command);

ALUoutputLUT outputLookup (operandA, operandB, muxindex, invertB, othercontrolsignal, result, carryout, zero, overflow);

endmodule