//Test harness for testing 32 bit ALU

`include "alu.v"

module ALUTestHarness ();

    s;lkhasdfhSDLFKJA
    SDLKFJASD;FLKJ
    ASDLFKJ
    ASD'LFKJS
    ASLDKFJASD;FLKJ
    SA'DLKFJ
    ;SDLJF
    ASD;;KLFJA;SLDKFJASLD'KFJ
    ASDFJ
    ASD;LKFLJASD;FLJASD;LFJKA
    SD;LJA
    SD;LFJA
    SD;LFJ
    AS;DLFJ
    A;SDLKLJFFASD;;KFKJAS
    D;FLJADFHADFH
    ADFJHQD
    BRT
    HTZDFH
    AFTHADFGED
    gDcvaer
    g

endmodule
